module alu(data_operandA, data_operandB, ctrl_ALUopcode, ctrl_shiftamt, data_result, isNotEqual, isLessThan, overflow);
        
    input [31:0] data_operandA, data_operandB;
    input [4:0] ctrl_ALUopcode, ctrl_shiftamt;

    output [31:0] data_result;
    output isNotEqual, isLessThan, overflow;

    // add your code here:
    
    wire [31:0] andresult;
    and and0(andresult[0], data_operandA[0], data_operandB[0]);
    and and1(andresult[1], data_operandA[1], data_operandB[1]);
    and and2(andresult[2], data_operandA[2], data_operandB[2]);
    and and3(andresult[3], data_operandA[3], data_operandB[3]);
    and and4(andresult[4], data_operandA[4], data_operandB[4]);
    and and5(andresult[5], data_operandA[5], data_operandB[5]);
    and and6(andresult[6], data_operandA[6], data_operandB[6]);
    and and7(andresult[7], data_operandA[7], data_operandB[7]);
    and and8(andresult[8], data_operandA[8], data_operandB[8]);
    and and9(andresult[9], data_operandA[9], data_operandB[9]);
    and and10(andresult[10], data_operandA[10], data_operandB[10]);
    and and11(andresult[11], data_operandA[11], data_operandB[11]);
    and and12(andresult[12], data_operandA[12], data_operandB[12]);
    and and13(andresult[13], data_operandA[13], data_operandB[13]);
    and and14(andresult[14], data_operandA[14], data_operandB[14]);
    and and15(andresult[15], data_operandA[15], data_operandB[15]);
    and and16(andresult[16], data_operandA[16], data_operandB[16]);
    and and17(andresult[17], data_operandA[17], data_operandB[17]);
    and and18(andresult[18], data_operandA[18], data_operandB[18]);
    and and19(andresult[19], data_operandA[19], data_operandB[19]);
    and and20(andresult[20], data_operandA[20], data_operandB[20]);
    and and21(andresult[21], data_operandA[21], data_operandB[21]);
    and and22(andresult[22], data_operandA[22], data_operandB[22]);
    and and23(andresult[23], data_operandA[23], data_operandB[23]);
    and and24(andresult[24], data_operandA[24], data_operandB[24]);
    and and25(andresult[25], data_operandA[25], data_operandB[25]);
    and and26(andresult[26], data_operandA[26], data_operandB[26]);
    and and27(andresult[27], data_operandA[27], data_operandB[27]);
    and and28(andresult[28], data_operandA[28], data_operandB[28]);
    and and29(andresult[29], data_operandA[29], data_operandB[29]);
    and and30(andresult[30], data_operandA[30], data_operandB[30]);
    and and31(andresult[31], data_operandA[31], data_operandB[31]);

    wire [31:0] orresult; 

    or or0(orresult[0], data_operandA[0], data_operandB[0]);
    or or1(orresult[1], data_operandA[1], data_operandB[1]);
    or or2(orresult[2], data_operandA[2], data_operandB[2]);
    or or3(orresult[3], data_operandA[3], data_operandB[3]);
    or or4(orresult[4], data_operandA[4], data_operandB[4]);
    or or5(orresult[5], data_operandA[5], data_operandB[5]);
    or or6(orresult[6], data_operandA[6], data_operandB[6]);
    or or7(orresult[7], data_operandA[7], data_operandB[7]);
    or or8(orresult[8], data_operandA[8], data_operandB[8]);
    or or9(orresult[9], data_operandA[9], data_operandB[9]);
    or or10(orresult[10], data_operandA[10], data_operandB[10]);
    or or11(orresult[11], data_operandA[11], data_operandB[11]);
    or or12(orresult[12], data_operandA[12], data_operandB[12]);
    or or13(orresult[13], data_operandA[13], data_operandB[13]);
    or or14(orresult[14], data_operandA[14], data_operandB[14]);
    or or15(orresult[15], data_operandA[15], data_operandB[15]);
    or or16(orresult[16], data_operandA[16], data_operandB[16]);
    or or17(orresult[17], data_operandA[17], data_operandB[17]);
    or or18(orresult[18], data_operandA[18], data_operandB[18]);
    or or19(orresult[19], data_operandA[19], data_operandB[19]);
    or or20(orresult[20], data_operandA[20], data_operandB[20]);
    or or21(orresult[21], data_operandA[21], data_operandB[21]);
    or or22(orresult[22], data_operandA[22], data_operandB[22]);
    or or23(orresult[23], data_operandA[23], data_operandB[23]);
    or or24(orresult[24], data_operandA[24], data_operandB[24]);
    or or25(orresult[25], data_operandA[25], data_operandB[25]);
    or or26(orresult[26], data_operandA[26], data_operandB[26]);
    or or27(orresult[27], data_operandA[27], data_operandB[27]);
    or or28(orresult[28], data_operandA[28], data_operandB[28]);
    or or29(orresult[29], data_operandA[29], data_operandB[29]);
    or or30(orresult[30], data_operandA[30], data_operandB[30]);
    or or31(orresult[31], data_operandA[31], data_operandB[31]);
   
    wire [31:0] lshiftresult;
    wire [31:0] lshift16, lshift8, lshift4, lshift2, lshift1, l16out, l8out, l4out, l2out;
    assign lshift16[31:16]= data_operandA[15:0];
    assign lshift16[15:0]=0;
    assign lshift8[7:0]=0;
    assign lshift4[3:0]=0;
    assign lshift2[1:0]=0;
    assign lshift1[0]=0;
    mux_2 l16(l16out, ctrl_shiftamt[4], data_operandA, lshift16);
    assign lshift8[31:8]= l16out[23:0];
    mux_2 l8(l8out, ctrl_shiftamt[3], l16out, lshift8);
    assign lshift4[31:4]= l8out[27:0];
    mux_2 l4(l4out, ctrl_shiftamt[2], l8out, lshift4);
    assign lshift2[31:2]= l4out[29:0];
    mux_2 l2(l2out, ctrl_shiftamt[1], l4out, lshift2);
    assign lshift1[31:1]= l2out[30:0];
    mux_2 l1(lshiftresult, ctrl_shiftamt[0], l2out, lshift1);
    wire [31:0] rshiftresult;
    wire [31:0] rshift16, rshift8, rshift4, rshift2, rshift1, r16out, r8out, r4out, r2out;
    assign rshift16[15:0]= data_operandA[31:16];
    assign rshift16[31]=data_operandA[31];
    assign rshift16[30]=data_operandA[31];
    assign rshift16[29]=data_operandA[31];
    assign rshift16[28]=data_operandA[31];
    assign rshift16[27]=data_operandA[31];
    assign rshift16[26]=data_operandA[31];
    assign rshift16[25]=data_operandA[31];
    assign rshift16[24]=data_operandA[31];
    assign rshift16[23]=data_operandA[31];
    assign rshift16[22]=data_operandA[31];
    assign rshift16[21]=data_operandA[31];
    assign rshift16[20]=data_operandA[31];
    assign rshift16[19]=data_operandA[31];
    assign rshift16[18]=data_operandA[31];
    assign rshift16[17]=data_operandA[31];
    assign rshift16[16]=data_operandA[31];
    assign rshift8[31]=data_operandA[31];
    assign rshift8[30]=data_operandA[31];
    assign rshift8[29]=data_operandA[31];
    assign rshift8[28]=data_operandA[31];
    assign rshift8[27]=data_operandA[31];
    assign rshift8[26]=data_operandA[31];
    assign rshift8[25]=data_operandA[31];
    assign rshift8[24]=data_operandA[31];
    assign rshift4[31]=data_operandA[31];
    assign rshift4[30]=data_operandA[31];
    assign rshift4[29]=data_operandA[31];
    assign rshift4[28]=data_operandA[31];
    assign rshift2[31]=data_operandA[31];
    assign rshift2[30]=data_operandA[31];
    assign rshift1[31]=data_operandA[31];
    mux_2 r16(r16out, ctrl_shiftamt[4], data_operandA, rshift16);
    assign rshift8[23:0]= r16out[31:8];
    mux_2 r8(r8out, ctrl_shiftamt[3], r16out, rshift8);
    assign rshift4[27:0]= r8out[31:4];
    mux_2 r4(r4out, ctrl_shiftamt[2], r8out, rshift4);
    assign rshift2[29:0]= r4out[31:2];
    mux_2 r2(r2out, ctrl_shiftamt[1], r4out, rshift2);
    assign rshift1[30:0]= r2out[31:1];
    mux_2 r1(rshiftresult, ctrl_shiftamt[0], r2out, rshift1);

    wire [31:0] addresult;
    wire carryzero, carryone, carrytwo, carrythree, carryfour;
    assign carryzero=0;
    eightbitCLA eight(addresult[7:0], carryone, data_operandA[7:0], data_operandB[7:0], carryzero);
    eightbitCLA sixteen(addresult[15:8], carrytwo, data_operandA[15:8], data_operandB[15:8], carryone);
    eightbitCLA twentyfour(addresult[23:16], carrythree, data_operandA[23:16], data_operandB[23:16], carrytwo);
    eightbitCLA thirtytwo(addresult[31:24], carryfour, data_operandA[31:24], data_operandB[31:24], carrythree);

    wire [31:0] subtractresult;
    wire scarryone, scarrytwo, scarrythree, scarryfour, scarryzero;
    assign scarryzero =1;
    wire [31:0] notdata_operandB;
    not n0(notdata_operandB[0], data_operandB[0]);
    not n1(notdata_operandB[1], data_operandB[1]);
    not n2(notdata_operandB[2], data_operandB[2]);
    not n3(notdata_operandB[3], data_operandB[3]);
    not n4(notdata_operandB[4], data_operandB[4]);
    not n5(notdata_operandB[5], data_operandB[5]);
    not n6(notdata_operandB[6], data_operandB[6]);
    not n7(notdata_operandB[7], data_operandB[7]);
    not n8(notdata_operandB[8], data_operandB[8]);
    not n9(notdata_operandB[9], data_operandB[9]);
    not n10(notdata_operandB[10], data_operandB[10]);
    not n11(notdata_operandB[11], data_operandB[11]);
    not n12(notdata_operandB[12], data_operandB[12]);
    not n13(notdata_operandB[13], data_operandB[13]);
    not n14(notdata_operandB[14], data_operandB[14]);
    not n15(notdata_operandB[15], data_operandB[15]);
    not n16(notdata_operandB[16], data_operandB[16]);
    not n17(notdata_operandB[17], data_operandB[17]);
    not n18(notdata_operandB[18], data_operandB[18]);
    not n19(notdata_operandB[19], data_operandB[19]);
    not n20(notdata_operandB[20], data_operandB[20]);
    not n21(notdata_operandB[21], data_operandB[21]);
    not n22(notdata_operandB[22], data_operandB[22]);
    not n23(notdata_operandB[23], data_operandB[23]);
    not n24(notdata_operandB[24], data_operandB[24]);
    not n25(notdata_operandB[25], data_operandB[25]);
    not n26(notdata_operandB[26], data_operandB[26]);
    not n27(notdata_operandB[27], data_operandB[27]);
    not n28(notdata_operandB[28], data_operandB[28]);
    not n29(notdata_operandB[29], data_operandB[29]);
    not n30(notdata_operandB[30], data_operandB[30]);
    not n31(notdata_operandB[31], data_operandB[31]);
   

    eightbitCLA seight(subtractresult[7:0], scarryone, data_operandA[7:0], notdata_operandB[7:0], scarryzero);
    eightbitCLA ssixteen(subtractresult[15:8], scarrytwo, data_operandA[15:8], notdata_operandB[15:8], scarryone);
    eightbitCLA stwentyfour(subtractresult[23:16], scarrythree, data_operandA[23:16], notdata_operandB[23:16], scarrytwo);
    eightbitCLA sthirtytwo(subtractresult[31:24], scarryfour, data_operandA[31:24], notdata_operandB[31:24], scarrythree);
     wire addoverflow, suboverflow, same, notsame, diff, secsame;
    mux_8 alumux(data_result, ctrl_ALUopcode[2:0], addresult, subtractresult, andresult, orresult, lshiftresult, rshiftresult, andresult, andresult);
    or noteq(isNotEqual, subtractresult[0], subtractresult[1], subtractresult[2], subtractresult[3], subtractresult[4], subtractresult[5], subtractresult[6], subtractresult[7], subtractresult[8], subtractresult[9], subtractresult[10], subtractresult[11], subtractresult[12], subtractresult[13], subtractresult[14], subtractresult[15], subtractresult[16], subtractresult[17], subtractresult[18], subtractresult[19], subtractresult[20], subtractresult[21], subtractresult[22], subtractresult[23], subtractresult[24], subtractresult[25], subtractresult[26], subtractresult[27], subtractresult[28], subtractresult[29], subtractresult[30], subtractresult[31]);
   
    xor diffsign(diff, data_operandA[31], data_operandB[31]);
    xnor samesign(same, data_operandA[31], data_operandB[31]);
    xor nsign(notsame, data_operandA[31], addresult[31]);
    and aover(addoverflow, notsame, same);
    xnor secsame(secsame, data_operandB[31], subtractresult[31]);
    and sover(suboverflow, secsame, diff);
    twomux_2 oselect(overflow, ctrl_ALUopcode[0], addoverflow, suboverflow);
    wire notover, check, bneg, notneg; 
    not nover(notover, overflow);
    and subcheck(check, subtractresult[31], notover);
    not aneg(notneg, data_operandB[31]);
    and bneg(bneg, notneg, data_operandA[31]);
    or less(isLessThan, check, bneg);
    
    


endmodule