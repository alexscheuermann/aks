module eightbitCLA(Sum, Carryout, A,B, Carryin);
    input [7:0] A, B;
    input Carryin; 
    output [7:0] Sum;
    output Carryout; 
    wire p7g6, p7p6g5, p7p6p5g4, p7p6p5p4g3, p7p6p5p4p3g2, p7p6p5p4p3p2g1, p7p6p5p4p3p2p1g0, p7p6p5p4p3p2p1p0c0, p6g5, p6p5g4, p6p5p4g3, p6p5p4p3g2, p6p5p4p3p2g1, p6p5p4p3p2p1g0, p6p5p4p3p2p1p0c0, p5g4, p5p4g3, p5p4p3g2, p5p4p3p2g1, p5p4p3p2p1g0, p5p4p3p2p1p0c0, p4g3, p4p3g2, p4p3p2g1, p4p3p2p1g0, p4p3p2p1p0c0, p3g2, p3p2g1, p3p2p1g0, p3p2p1p0c0, p2g1, p2p1g0, p2p1p0c0, p1p0c0, p1g0, p0c0, g0, p0, c1, c2, c3, c4, c5, c6, c7, g1, p1, g2, p2, g3, p3, g4, p4, g5, p5, g6, p6, g7, p7; 
    and gen0(g0, A[0], B[0]);
    or prop0(p0, A[0], B[0]);
    and gen1(g1, A[1], B[1]);
    or prop1(p1, A[1], B[1]);
    and gen2(g2, A[2], B[2]);
    or prop2(p2, A[2], B[2]);
    and gen3(g3, A[3], B[3]);
    or prop3(p3, A[3], B[3]);
    and gen4(g4, A[4], B[4]);
    or prop4(p4, A[4], B[4]);
    and gen5(g5, A[5], B[5]);
    or prop5(p5, A[5], B[5]);
    and gen6(g6, A[6], B[6]);
    or prop6(p6, A[6], B[6]);
    and gen7(g7, A[7], B[7]);
    or prop7(p7, A[7], B[7]);
    and p0c0(p0c0, p0, Carryin);
    or c1(c1, p0c0,g0);
    and p1g0(p1g0, p1, g0);
    and p1p0c0(p1p0c0, p1, p0, Carryin);
    or c2(c2, g1, p1g0, p1p0c0);
    and p2g1 (p2g1, p2, g1);
    and p2p1g0(p2p1g0, p2, p1, g0);
    and p2p1p0c0(p2p1p0c0, p2, p1, p0, Carryin);
    or c3(c3, g2, p2g1, p2p1g0,p2p1p0c0);
    and p3g2(p3g2, p3, g2);
    and p3p2g1 (p3p2g1, p3, p2, g1);
    and p3p2p1g0(p3p2p1g0, p3, p2, p1, g0);
    and p3p2p1p0c0(p3p2p1p0c0, p3, p2, p1, p0, Carryin);
    or c4(c4, g3, p3g2, p3p2g1, p3p2p1g0, p3p2p1p0c0);
    and p4g3 (p4g3, p4, g3);
    and p4p3g2 (p4p3g2, p4, p3, g2);
    and p4p3p2g1(p4p3p2g1, p4, p3, p2, g1);
    and p4p3p2p1g0(p4p3p2p1g0, p4, p3, p2, p1, g0);
    and p4p3p2p1p0c0(p4p3p2p1p0c0, p4, p3, p2, p1, p0, Carryin);
    or  c5(c5, g4, p4g3, p4p3g2, p4p3p2g1, p4p3p2p1g0, p4p3p2p1p0c0);
    and p5g4 (p5g4, p5, g4);
    and p5p4g3 (p5p4g3, p5, p4, g3);
    and p5p4p3g2 (p5p4p3g2, p5, p4, p3, g2);
    and p5p4p3p2g1(p5p4p3p2g1, p5, p4, p3, p2, g1);
    and p5p4p3p2p1g0(p5p4p3p2p1g0, p5, p4, p3, p2, p1, g0);
    and p5p4p3p2p1p0c0(p5p4p3p2p1p0c0, p5, p4, p3, p2, p1, p0, Carryin);
    or  c6(c6, g5, p5g4, p5p4g3, p5p4p3g2, p5p4p3p2g1, p5p4p3p2p1g0, p5p4p3p2p1p0c0);
    and p6g5 (p6g5, p6, g5);
    and p6p5g4 (p6p5g4, p6, p5, g4);
    and p6p5p4g3 (p6p5p4g3, p6, p5, p4, g3);
    and p6p5p4p3g2 (p6p5p4p3g2, p6, p5, p4, p3, g2);
    and p6p5p4p3p2g1(p6p5p4p3p2g1, p6, p5, p4, p3, p2, g1);
    and p6p5p4p3p2p1g0(p6p5p4p3p2p1g0, p6, p5, p4, p3, p2, p1, g0);
    and p6p5p4p3p2p1p0c0(p6p5p4p3p2p1p0c0, p6, p5, p4, p3, p2, p1, p0, Carryin);
    or  c7(c7, g6, p6g5, p6p5g4, p6p5p4g3, p6p5p4p3g2, p6p5p4p3p2g1, p6p5p4p3p2p1g0, p6p5p4p3p2p1p0c0);
    and p7g6 (p7g6, p7, g6);
    and p7p6g5 (p7p6g5, p7, p6, g5);
    and p7p6p5g4 (p7p6p5g4, p7, p6, p5, g4);
    and p7p6p5p4g3 (p7p6p5p4g3, p7, p6, p5, p4, g3);
    and p7p6p5p4p3g2 (p7p6p5p4p3g2, p7, p6, p5, p4, p3, g2);
    and p7p6p5p4p3p2g1(p7p6p5p4p3p2g1, p7, p6, p5, p4, p3, p2, g1);
    and p7p6p5p4p3p2p1g0(p7p6p5p4p3p2p1g0, p7, p6, p5, p4, p3, p2, p1, g0);
    and p7p6p5p4p3p2p1p0c0(p7p6p5p4p3p2p1p0c0, p7, p6, p5, p4, p3, p2, p1, p0, Carryin);
    or  cout(Carryout, g7, p7g6, p7p6g5, p7p6p5g4, p7p6p5p4g3, p7p6p5p4p3g2, p7p6p5p4p3p2g1, p7p6p5p4p3p2p1g0, p7p6p5p4p3p2p1p0c0);
    xor sum0(Sum[0], Carryin, A[0], B[0]);
    xor sum1(Sum[1], c1, A[1], B[1]);
    xor sum2(Sum[2], c2, A[2], B[2]);
    xor sum3(Sum[3], c3, A[3], B[3]);
    xor sum4(Sum[4], c4, A[4], B[4]);
    xor sum5(Sum[5], c5, A[5], B[5]);
    xor sum6(Sum[6], c6, A[6], B[6]);
    xor sum7(Sum[7], c7, A[7], B[7]);
endmodule